module memory(clk,
              rst,
              aw_id
              );

end module
