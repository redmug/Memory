module 

end module

